library verilog;
use verilog.vl_types.all;
entity csb_vlg_vec_tst is
end csb_vlg_vec_tst;
